library ieee;
use ieee.std_logic_1164.all;

entity detector is
port( x: in std_logic_vector(3 downto 0);
		y: out std_logic_vector(0 downto 0));

end detector;

architecture a1 of detector is
begin
detector: process(x)
begin
if x = "0000" then 
	y <= "1";
elsif x = "0100" then
	y <= "1";
elsif x = "1000" then 
   y <= "1";
elsif x = "1110" then 
   y <= "1";	
else y <= "0";
end if;
end process;
end a1;
